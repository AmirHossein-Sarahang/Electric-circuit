** Profile: "SCHEMATIC1-soal5"  [ C:\USERS\ARIAN 3\DESKTOP\PROJE1\5\soal5-SCHEMATIC1-soal5.sim ] 

** Creating circuit file "soal5-SCHEMATIC1-soal5.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 2000 1 10000k
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\soal5-SCHEMATIC1.net" 


.END
