** Profile: "SCHEMATIC1-soal1"  [ C:\Users\arian 3\Desktop\proje1\soal1-SCHEMATIC1-soal1.sim ] 

** Creating circuit file "soal1-SCHEMATIC1-soal1.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 100ms 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\soal1-SCHEMATIC1.net" 


.END
