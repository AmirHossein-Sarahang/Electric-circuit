** Profile: "SCHEMATIC1-soal3"  [ C:\USERS\ARIAN 3\DESKTOP\PROJE1\3\soal3-SCHEMATIC1-soal3.sim ] 

** Creating circuit file "soal3-SCHEMATIC1-soal3.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 2000 1 100000k
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\soal3-SCHEMATIC1.net" 


.END
