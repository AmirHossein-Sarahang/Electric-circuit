** Profile: "SCHEMATIC1-soal6"  [ C:\USERS\ARIAN 3\DESKTOP\PROJE1\6\soal6-SCHEMATIC1-soal6.sim ] 

** Creating circuit file "soal6-SCHEMATIC1-soal6.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 2000 1 10000k
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\soal6-SCHEMATIC1.net" 


.END
