** Profile: "SCHEMATIC1-soal4"  [ C:\USERS\ARIAN 3\DESKTOP\PROJE1\4\soal4-SCHEMATIC1-soal4.sim ] 

** Creating circuit file "soal4-SCHEMATIC1-soal4.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC DEC PARAM Rvar 1 10k 20 
+ DEC PARAM Rvar1 1 10k 20 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\soal4-SCHEMATIC1.net" 


.END
